* 2-input NAND gate
.title CMOS NAND Gate

.param vdd=1.8

* Inputs
Vin1 a 0 PULSE(0 {vdd} 0ns 0.1ns 0.1ns 10ns 20ns)
Vin2 b 0 PULSE(0 {vdd} 0ns 0.1ns 0.1ns 20ns 40ns)

* PMOS transistors (parallel - pull-up network)
M1 out a vdd vdd pmos W=2u L=180n
M2 out b vdd vdd pmos W=2u L=180n

* NMOS transistors (series - pull-down network)
M3 out a n1 0 nmos W=1u L=180n
M4 n1 b 0 0 nmos W=1u L=180n

* Load
Cload out 0 10fF
Vdd vdd 0 DC {vdd}

.model nmos NMOS (Level=1 VTO=0.4 KP=120u)
.model pmos PMOS (Level=1 VTO=-0.4 KP=40u)

.tran 0.01ns 80ns
.control
run
plot v(a) v(b) v(out)
.endc
.end

